module regfile_tb();
		logic clk,we3;
		logic [4:0] ra1,ra2,wa3;
		logic [63:0] wd3, rd1, rd2;
		
	
	regfile dut(clk, we3, ra1, ra2, wa3, wd3, rd1, rd2);
	//clock generation @100MHz 10ns
	always
		begin
				clk = 1; #10; clk=0; #10;
		end
	
	initial