module maindec_tb();

endmodule