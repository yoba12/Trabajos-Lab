module allu_tb();

endmodule